

module A2DFFQN_X0P5M (A, B, CK, QN);

	//ports
	input A;
	input B;
	input CK;
	output QN;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;

endmodule


module A2DFFQN_X1M (A, B, CK, QN);

	//ports
	input A;
	input B;
	input CK;
	output QN;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;

endmodule


module A2DFFQN_X2M (A, B, CK, QN);

	//ports
	input A;
	input B;
	input CK;
	output QN;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;

endmodule


module A2DFFQN_X3M (A, B, CK, QN);

	//ports
	input A;
	input B;
	input CK;
	output QN;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;

endmodule


module A2DFFQ_X0P5M (A, B, CK, Q);

	//ports
	input A;
	input B;
	input CK;
	output Q;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;

endmodule


module A2DFFQ_X1M (A, B, CK, Q);

	//ports
	input A;
	input B;
	input CK;
	output Q;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;

endmodule


module A2DFFQ_X2M (A, B, CK, Q);

	//ports
	input A;
	input B;
	input CK;
	output Q;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;

endmodule


module A2DFFQ_X3M (A, B, CK, Q);

	//ports
	input A;
	input B;
	input CK;
	output Q;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;

endmodule


module A2DFFQ_X4M (A, B, CK, Q);

	//ports
	input A;
	input B;
	input CK;
	output Q;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;

endmodule


module A2SDFFQN_X0P5M (A, B, CK, QN, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output QN;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;
	wire SE;
	wire SI;

endmodule


module A2SDFFQN_X1M (A, B, CK, QN, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output QN;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;
	wire SE;
	wire SI;

endmodule


module A2SDFFQN_X2M (A, B, CK, QN, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output QN;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;
	wire SE;
	wire SI;

endmodule


module A2SDFFQN_X3M (A, B, CK, QN, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output QN;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire QN;
	wire SE;
	wire SI;

endmodule


module A2SDFFQ_X0P5M (A, B, CK, Q, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output Q;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;
	wire SE;
	wire SI;

endmodule


module A2SDFFQ_X1M (A, B, CK, Q, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output Q;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;
	wire SE;
	wire SI;

endmodule


module A2SDFFQ_X2M (A, B, CK, Q, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output Q;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;
	wire SE;
	wire SI;

endmodule


module A2SDFFQ_X3M (A, B, CK, Q, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output Q;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;
	wire SE;
	wire SI;

endmodule


module A2SDFFQ_X4M (A, B, CK, Q, SE, SI);

	//ports
	input A;
	input B;
	input CK;
	output Q;
	input SE;
	input SI;

	//wires
	wire A;
	wire B;
	wire CK;
	wire Q;
	wire SE;
	wire SI;

endmodule


module ADDFCIN_X1M (A, B, CIN, CO, SUM);

	//ports
	input A;
	input B;
	input CIN;
	output CO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire CIN;
	wire CO;
	wire SUM;

endmodule


module ADDFCIN_X1P4M (A, B, CIN, CO, SUM);

	//ports
	input A;
	input B;
	input CIN;
	output CO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire CIN;
	wire CO;
	wire SUM;

endmodule


module ADDFCIN_X2M (A, B, CIN, CO, SUM);

	//ports
	input A;
	input B;
	input CIN;
	output CO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire CIN;
	wire CO;
	wire SUM;

endmodule


module ADDFH_X1M (A, B, CI, CO, SUM);

	//ports
	input A;
	input B;
	input CI;
	output CO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;
	wire SUM;

endmodule


module ADDFH_X1P4M (A, B, CI, CO, SUM);

	//ports
	input A;
	input B;
	input CI;
	output CO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;
	wire SUM;

endmodule


module ADDFH_X2M (A, B, CI, CO, SUM);

	//ports
	input A;
	input B;
	input CI;
	output CO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;
	wire SUM;

endmodule


module ADDF_X1M (A, B, CI, CO, S);

	//ports
	input A;
	input B;
	input CI;
	output CO;
	output S;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;
	wire S;

endmodule


module ADDF_X1P4M (A, B, CI, CO, S);

	//ports
	input A;
	input B;
	input CI;
	output CO;
	output S;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;
	wire S;

endmodule


module ADDF_X2M (A, B, CI, CO, S);

	//ports
	input A;
	input B;
	input CI;
	output CO;
	output S;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;
	wire S;

endmodule


module ADDH_X1M (A, B, CO, S);

	//ports
	input A;
	input B;
	output CO;
	output S;

	//wires
	wire A;
	wire B;
	wire CO;
	wire S;

endmodule


module ADDH_X1P4M (A, B, CO, S);

	//ports
	input A;
	input B;
	output CO;
	output S;

	//wires
	wire A;
	wire B;
	wire CO;
	wire S;

endmodule


module ADDH_X2M (A, B, CO, S);

	//ports
	input A;
	input B;
	output CO;
	output S;

	//wires
	wire A;
	wire B;
	wire CO;
	wire S;

endmodule


module AND2_X0P5M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X0P7M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X11M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X1M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X1P4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X2M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X3M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X6M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND2_X8M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module AND3_X0P5M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X0P7M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X11M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X1M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X1P4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X2M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X3M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X6M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND3_X8M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module AND4_X0P5M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X0P7M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X1M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X1P4M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X2M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X3M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X4M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X6M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module AND4_X8M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module ANTENNA2 (A);

	//ports
	input A;

	//wires
	wire A;

endmodule


module AO1B2_X0P5M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X0P7M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X1M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X1P4M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X2M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X3M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X4M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO1B2_X6M (A0N, B0, B1, Y);

	//ports
	input A0N;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0N;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO21B_X0P5M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X0P7M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X1M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X1P4M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X2M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X3M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X4M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21B_X6M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AO21_X0P5M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X0P7M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X1M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X1P4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X2M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X3M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO21_X6M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AO22_X0P5M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X0P7M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X1M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X1P4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X2M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X3M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AO22_X6M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI211_X0P5M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI211_X0P7M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI211_X1M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI211_X1P4M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI211_X2M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI211_X3M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI211_X4M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module AOI21B_X0P5M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X0P7M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X1M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X1P4M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X2M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X3M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X4M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X6M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21B_X8M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module AOI21_X0P5M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X0P7M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X1M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X1P4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X2M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X3M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X6M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI21_X8M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module AOI221_X0P5M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI221_X0P7M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI221_X1M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI221_X1P4M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI221_X2M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI221_X3M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI221_X4M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module AOI222_X0P5M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI222_X0P7M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI222_X1M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI222_X1P4M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI222_X2M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI222_X3M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI222_X4M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module AOI22_X0P5M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X0P7M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X1M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X1P4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X2M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X3M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X6M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI22_X8M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI2XB1_X0P5M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X0P7M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X1M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X1P4M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X2M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X3M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X4M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X6M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI2XB1_X8M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module AOI31_X0P5M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X0P7M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X1M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X1P4M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X2M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X3M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X4M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI31_X6M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module AOI32_X0P5M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X0P7M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X1M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X1P4M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X2M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X3M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X4M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module AOI32_X6M (A0, A1, A2, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire B1;
	wire Y;

endmodule


module BENC_X11M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BENC_X16M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BENC_X2M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BENC_X3M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BENC_X4M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BENC_X6M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BENC_X8M (AN, M0, M1, M2, SN, X2);

	//ports
	output AN;
	input M0;
	input M1;
	input M2;
	output SN;
	output X2;

	//wires
	wire AN;
	wire M0;
	wire M1;
	wire M2;
	wire SN;
	wire X2;

endmodule


module BMXIT_X0P7M (AN, D0, D1, PPN, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PPN;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PPN;
	wire SN;
	wire X2;

endmodule


module BMXIT_X1M (AN, D0, D1, PPN, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PPN;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PPN;
	wire SN;
	wire X2;

endmodule


module BMXIT_X1P4M (AN, D0, D1, PPN, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PPN;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PPN;
	wire SN;
	wire X2;

endmodule


module BMXIT_X2M (AN, D0, D1, PPN, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PPN;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PPN;
	wire SN;
	wire X2;

endmodule


module BMXT_X0P7M (AN, D0, D1, PP, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PP;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PP;
	wire SN;
	wire X2;

endmodule


module BMXT_X1M (AN, D0, D1, PP, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PP;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PP;
	wire SN;
	wire X2;

endmodule


module BMXT_X1P4M (AN, D0, D1, PP, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PP;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PP;
	wire SN;
	wire X2;

endmodule


module BMXT_X2M (AN, D0, D1, PP, SN, X2);

	//ports
	input AN;
	input D0;
	input D1;
	output PP;
	input SN;
	input X2;

	//wires
	wire AN;
	wire D0;
	wire D1;
	wire PP;
	wire SN;
	wire X2;

endmodule


module BUFH_X0P7M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X0P8M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X11M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X13M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X16M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X1M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X1P2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X1P4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X1P7M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X2P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X3M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X3P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X6M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X7P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFH_X9M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUFZ_X11M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X16M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X1M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X1P4M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X2M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X3M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X4M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X6M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUFZ_X8M (A, OE, Y);

	//ports
	input A;
	input OE;
	output Y;

	//wires
	wire A;
	wire OE;
	wire Y;

endmodule


module BUF_X0P7B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X0P7M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X0P8B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X0P8M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X11B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X11M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X13B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X13M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X16B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X16M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1P2B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1P2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1P4B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1P4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1P7B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X1P7M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X2B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X2P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X2P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X3B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X3M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X3P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X3P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X4B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X6B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X6M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X7P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X7P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X9B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module BUF_X9M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module CGENCIN_X1M (A, B, CIN, CO);

	//ports
	input A;
	input B;
	input CIN;
	output CO;

	//wires
	wire A;
	wire B;
	wire CIN;
	wire CO;

endmodule


module CGENCIN_X1P4M (A, B, CIN, CO);

	//ports
	input A;
	input B;
	input CIN;
	output CO;

	//wires
	wire A;
	wire B;
	wire CIN;
	wire CO;

endmodule


module CGENCIN_X2M (A, B, CIN, CO);

	//ports
	input A;
	input B;
	input CIN;
	output CO;

	//wires
	wire A;
	wire B;
	wire CIN;
	wire CO;

endmodule


module CGENCON_X1M (A, B, CI, CON);

	//ports
	input A;
	input B;
	input CI;
	output CON;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CON;

endmodule


module CGENCON_X1P4M (A, B, CI, CON);

	//ports
	input A;
	input B;
	input CI;
	output CON;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CON;

endmodule


module CGENCON_X2M (A, B, CI, CON);

	//ports
	input A;
	input B;
	input CI;
	output CON;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CON;

endmodule


module CGENI_X1M (A, B, CI, CON);

	//ports
	input A;
	input B;
	input CI;
	output CON;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CON;

endmodule


module CGENI_X1P4M (A, B, CI, CON);

	//ports
	input A;
	input B;
	input CI;
	output CON;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CON;

endmodule


module CGENI_X2M (A, B, CI, CON);

	//ports
	input A;
	input B;
	input CI;
	output CON;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CON;

endmodule


module CGEN_X1M (A, B, CI, CO);

	//ports
	input A;
	input B;
	input CI;
	output CO;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;

endmodule


module CGEN_X1P4M (A, B, CI, CO);

	//ports
	input A;
	input B;
	input CI;
	output CO;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;

endmodule


module CGEN_X2M (A, B, CI, CO);

	//ports
	input A;
	input B;
	input CI;
	output CO;

	//wires
	wire A;
	wire B;
	wire CI;
	wire CO;

endmodule


module CMPR42_X1M (A, B, C, CO, D, ICI, ICO, SUM);

	//ports
	input A;
	input B;
	input C;
	output CO;
	input D;
	input ICI;
	output ICO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire C;
	wire CO;
	wire D;
	wire ICI;
	wire ICO;
	wire SUM;

endmodule


module CMPR42_X1P4M (A, B, C, CO, D, ICI, ICO, SUM);

	//ports
	input A;
	input B;
	input C;
	output CO;
	input D;
	input ICI;
	output ICO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire C;
	wire CO;
	wire D;
	wire ICI;
	wire ICO;
	wire SUM;

endmodule


module CMPR42_X2M (A, B, C, CO, D, ICI, ICO, SUM);

	//ports
	input A;
	input B;
	input C;
	output CO;
	input D;
	input ICI;
	output ICO;
	output SUM;

	//wires
	wire A;
	wire B;
	wire C;
	wire CO;
	wire D;
	wire ICI;
	wire ICO;
	wire SUM;

endmodule


module DFFNQ_X1M (CKN, D, Q);

	//ports
	input CKN;
	input D;
	output Q;

	//wires
	wire CKN;
	wire D;
	wire Q;

endmodule


module DFFNQ_X2M (CKN, D, Q);

	//ports
	input CKN;
	input D;
	output Q;

	//wires
	wire CKN;
	wire D;
	wire Q;

endmodule


module DFFNQ_X3M (CKN, D, Q);

	//ports
	input CKN;
	input D;
	output Q;

	//wires
	wire CKN;
	wire D;
	wire Q;

endmodule


module DFFNRPQ_X1M (CKN, D, Q, R);

	//ports
	input CKN;
	input D;
	output Q;
	input R;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFNRPQ_X2M (CKN, D, Q, R);

	//ports
	input CKN;
	input D;
	output Q;
	input R;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFNRPQ_X3M (CKN, D, Q, R);

	//ports
	input CKN;
	input D;
	output Q;
	input R;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFNSQ_X1M (CKN, D, Q, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFNSQ_X2M (CKN, D, Q, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFNSQ_X3M (CKN, D, Q, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFNSRPQ_X1M (CKN, D, Q, R, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFNSRPQ_X2M (CKN, D, Q, R, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFNSRPQ_X3M (CKN, D, Q, R, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFQN_X0P5M (CK, D, QN);

	//ports
	input CK;
	input D;
	output QN;

	//wires
	wire CK;
	wire D;
	wire QN;

endmodule


module DFFQN_X1M (CK, D, QN);

	//ports
	input CK;
	input D;
	output QN;

	//wires
	wire CK;
	wire D;
	wire QN;

endmodule


module DFFQN_X2M (CK, D, QN);

	//ports
	input CK;
	input D;
	output QN;

	//wires
	wire CK;
	wire D;
	wire QN;

endmodule


module DFFQN_X3M (CK, D, QN);

	//ports
	input CK;
	input D;
	output QN;

	//wires
	wire CK;
	wire D;
	wire QN;

endmodule


module DFFQ_X0P5M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFQ_X1M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFQ_X2M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFQ_X3M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFQ_X4M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFRPQN_X0P5M (CK, D, QN, R);

	//ports
	input CK;
	input D;
	output QN;
	input R;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;

endmodule


module DFFRPQN_X1M (CK, D, QN, R);

	//ports
	input CK;
	input D;
	output QN;
	input R;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;

endmodule


module DFFRPQN_X2M (CK, D, QN, R);

	//ports
	input CK;
	input D;
	output QN;
	input R;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;

endmodule


module DFFRPQN_X3M (CK, D, QN, R);

	//ports
	input CK;
	input D;
	output QN;
	input R;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;

endmodule


module DFFRPQ_X0P5M (CK, D, Q, R);

	//ports
	input CK;
	input D;
	output Q;
	input R;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFRPQ_X1M (CK, D, Q, R);

	//ports
	input CK;
	input D;
	output Q;
	input R;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFRPQ_X2M (CK, D, Q, R);

	//ports
	input CK;
	input D;
	output Q;
	input R;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFRPQ_X3M (CK, D, Q, R);

	//ports
	input CK;
	input D;
	output Q;
	input R;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFRPQ_X4M (CK, D, Q, R);

	//ports
	input CK;
	input D;
	output Q;
	input R;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;

endmodule


module DFFSQN_X0P5M (CK, D, QN, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SN;

endmodule


module DFFSQN_X1M (CK, D, QN, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SN;

endmodule


module DFFSQN_X2M (CK, D, QN, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SN;

endmodule


module DFFSQN_X3M (CK, D, QN, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SN;

endmodule


module DFFSQ_X0P5M (CK, D, Q, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFSQ_X1M (CK, D, Q, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFSQ_X2M (CK, D, Q, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFSQ_X3M (CK, D, Q, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFSQ_X4M (CK, D, Q, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SN;

endmodule


module DFFSRPQ_X0P5M (CK, D, Q, R, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFSRPQ_X1M (CK, D, Q, R, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFSRPQ_X2M (CK, D, Q, R, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFSRPQ_X3M (CK, D, Q, R, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFSRPQ_X4M (CK, D, Q, R, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SN;

endmodule


module DFFYQ_X1M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFYQ_X2M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFYQ_X3M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DFFYQ_X4M (CK, D, Q);

	//ports
	input CK;
	input D;
	output Q;

	//wires
	wire CK;
	wire D;
	wire Q;

endmodule


module DLY2_X0P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY2_X1M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY2_X2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY2_X4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY4_X0P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY4_X1M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY4_X2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module DLY4_X4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module EDFFQN_X0P5M (CK, D, E, QN);

	//ports
	input CK;
	input D;
	input E;
	output QN;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;

endmodule


module EDFFQN_X1M (CK, D, E, QN);

	//ports
	input CK;
	input D;
	input E;
	output QN;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;

endmodule


module EDFFQN_X2M (CK, D, E, QN);

	//ports
	input CK;
	input D;
	input E;
	output QN;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;

endmodule


module EDFFQN_X3M (CK, D, E, QN);

	//ports
	input CK;
	input D;
	input E;
	output QN;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;

endmodule


module EDFFQ_X0P5M (CK, D, E, Q);

	//ports
	input CK;
	input D;
	input E;
	output Q;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;

endmodule


module EDFFQ_X1M (CK, D, E, Q);

	//ports
	input CK;
	input D;
	input E;
	output Q;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;

endmodule


module EDFFQ_X2M (CK, D, E, Q);

	//ports
	input CK;
	input D;
	input E;
	output Q;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;

endmodule


module EDFFQ_X3M (CK, D, E, Q);

	//ports
	input CK;
	input D;
	input E;
	output Q;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;

endmodule


module ENDCAPTIE2 ();

	//wires

endmodule


module ESDFFQN_X0P5M (CK, D, E, QN, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;
	wire SE;
	wire SI;

endmodule


module ESDFFQN_X1M (CK, D, E, QN, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;
	wire SE;
	wire SI;

endmodule


module ESDFFQN_X2M (CK, D, E, QN, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;
	wire SE;
	wire SI;

endmodule


module ESDFFQN_X3M (CK, D, E, QN, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire QN;
	wire SE;
	wire SI;

endmodule


module ESDFFQ_X0P5M (CK, D, E, Q, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;
	wire SE;
	wire SI;

endmodule


module ESDFFQ_X1M (CK, D, E, Q, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;
	wire SE;
	wire SI;

endmodule


module ESDFFQ_X2M (CK, D, E, Q, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;
	wire SE;
	wire SI;

endmodule


module ESDFFQ_X3M (CK, D, E, Q, SE, SI);

	//ports
	input CK;
	input D;
	input E;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire E;
	wire Q;
	wire SE;
	wire SI;

endmodule


module FILL128 ();

	//wires

endmodule


module FILL16 ();

	//wires

endmodule


module FILL1 ();

	//wires

endmodule


module FILL25CAP128 ();

	//wires

endmodule


module FILL25CAP12 ();

	//wires

endmodule


module FILL25CAP16 ();

	//wires

endmodule


module FILL25CAP32 ();

	//wires

endmodule


module FILL25CAP64 ();

	//wires

endmodule


module FILL25CAPTIE128 ();

	//wires

endmodule


module FILL25CAPTIE12 ();

	//wires

endmodule


module FILL25CAPTIE16 ();

	//wires

endmodule


module FILL25CAPTIE32 ();

	//wires

endmodule


module FILL25CAPTIE64 ();

	//wires

endmodule


module FILL2 ();

	//wires

endmodule


module FILL32 ();

	//wires

endmodule


module FILL4 ();

	//wires

endmodule


module FILL64 ();

	//wires

endmodule


module FILL8 ();

	//wires

endmodule


module FILLCAP128 ();

	//wires

endmodule


module FILLCAP16 ();

	//wires

endmodule


module FILLCAP32 ();

	//wires

endmodule


module FILLCAP3 ();

	//wires

endmodule


module FILLCAP4 ();

	//wires

endmodule


module FILLCAP64 ();

	//wires

endmodule


module FILLCAP8 ();

	//wires

endmodule


module FILLCAPTIE128 ();

	//wires

endmodule


module FILLCAPTIE16 ();

	//wires

endmodule


module FILLCAPTIE32 ();

	//wires

endmodule


module FILLCAPTIE64 ();

	//wires

endmodule


module FILLCAPTIE6 ();

	//wires

endmodule


module FILLCAPTIE8 ();

	//wires

endmodule


module FILLTIE128 ();

	//wires

endmodule


module FILLTIE16 ();

	//wires

endmodule


module FILLTIE2 ();

	//wires

endmodule


module FILLTIE32 ();

	//wires

endmodule


module FILLTIE4 ();

	//wires

endmodule


module FILLTIE64 ();

	//wires

endmodule


module FILLTIE8 ();

	//wires

endmodule


module FRICG_X0P5B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X0P6B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X0P7B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X0P8B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X11B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X13B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X16B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X1B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X1P2B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X1P4B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X1P7B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X2B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X2P5B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X3B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X3P5B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X4B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X5B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X6B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X7P5B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module FRICG_X9B (CK, ECK);

	//ports
	input CK;
	output ECK;

	//wires
	wire CK;
	wire ECK;

endmodule


module INV_X0P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P6B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P6M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P7B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P7M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P8B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X0P8M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X11B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X11M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X13B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X13M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X16B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X16M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1P2B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1P2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1P4B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1P4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1P7B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X1P7M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X2B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X2M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X2P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X2P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X3B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X3M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X3P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X3P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X4B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X4M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X6B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X6M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X7P5B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X7P5M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X9B (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module INV_X9M (A, Y);

	//ports
	input A;
	output Y;

	//wires
	wire A;
	wire Y;

endmodule


module LATNQN_X0P5M (D, GN, QN);

	//ports
	input D;
	input GN;
	output QN;

	//wires
	wire D;
	wire GN;
	wire QN;

endmodule


module LATNQN_X1M (D, GN, QN);

	//ports
	input D;
	input GN;
	output QN;

	//wires
	wire D;
	wire GN;
	wire QN;

endmodule


module LATNQN_X2M (D, GN, QN);

	//ports
	input D;
	input GN;
	output QN;

	//wires
	wire D;
	wire GN;
	wire QN;

endmodule


module LATNQN_X3M (D, GN, QN);

	//ports
	input D;
	input GN;
	output QN;

	//wires
	wire D;
	wire GN;
	wire QN;

endmodule


module LATNQN_X4M (D, GN, QN);

	//ports
	input D;
	input GN;
	output QN;

	//wires
	wire D;
	wire GN;
	wire QN;

endmodule


module LATNQ_X0P5M (D, GN, Q);

	//ports
	input D;
	input GN;
	output Q;

	//wires
	wire D;
	wire GN;
	wire Q;

endmodule


module LATNQ_X1M (D, GN, Q);

	//ports
	input D;
	input GN;
	output Q;

	//wires
	wire D;
	wire GN;
	wire Q;

endmodule


module LATNQ_X2M (D, GN, Q);

	//ports
	input D;
	input GN;
	output Q;

	//wires
	wire D;
	wire GN;
	wire Q;

endmodule


module LATNQ_X3M (D, GN, Q);

	//ports
	input D;
	input GN;
	output Q;

	//wires
	wire D;
	wire GN;
	wire Q;

endmodule


module LATNRPQN_X0P5M (D, GN, QN, R);

	//ports
	input D;
	input GN;
	output QN;
	input R;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire R;

endmodule


module LATNRPQN_X1M (D, GN, QN, R);

	//ports
	input D;
	input GN;
	output QN;
	input R;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire R;

endmodule


module LATNRPQN_X2M (D, GN, QN, R);

	//ports
	input D;
	input GN;
	output QN;
	input R;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire R;

endmodule


module LATNRPQN_X3M (D, GN, QN, R);

	//ports
	input D;
	input GN;
	output QN;
	input R;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire R;

endmodule


module LATNRPQN_X4M (D, GN, QN, R);

	//ports
	input D;
	input GN;
	output QN;
	input R;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire R;

endmodule


module LATNRQ_X0P5M (D, GN, Q, RN);

	//ports
	input D;
	input GN;
	output Q;
	input RN;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire RN;

endmodule


module LATNRQ_X1M (D, GN, Q, RN);

	//ports
	input D;
	input GN;
	output Q;
	input RN;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire RN;

endmodule


module LATNRQ_X2M (D, GN, Q, RN);

	//ports
	input D;
	input GN;
	output Q;
	input RN;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire RN;

endmodule


module LATNRQ_X3M (D, GN, Q, RN);

	//ports
	input D;
	input GN;
	output Q;
	input RN;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire RN;

endmodule


module LATNSPQ_X0P5M (D, GN, Q, S);

	//ports
	input D;
	input GN;
	output Q;
	input S;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire S;

endmodule


module LATNSPQ_X1M (D, GN, Q, S);

	//ports
	input D;
	input GN;
	output Q;
	input S;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire S;

endmodule


module LATNSPQ_X2M (D, GN, Q, S);

	//ports
	input D;
	input GN;
	output Q;
	input S;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire S;

endmodule


module LATNSPQ_X3M (D, GN, Q, S);

	//ports
	input D;
	input GN;
	output Q;
	input S;

	//wires
	wire D;
	wire GN;
	wire Q;
	wire S;

endmodule


module LATNSQN_X0P5M (D, GN, QN, SN);

	//ports
	input D;
	input GN;
	output QN;
	input SN;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire SN;

endmodule


module LATNSQN_X1M (D, GN, QN, SN);

	//ports
	input D;
	input GN;
	output QN;
	input SN;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire SN;

endmodule


module LATNSQN_X2M (D, GN, QN, SN);

	//ports
	input D;
	input GN;
	output QN;
	input SN;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire SN;

endmodule


module LATNSQN_X3M (D, GN, QN, SN);

	//ports
	input D;
	input GN;
	output QN;
	input SN;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire SN;

endmodule


module LATNSQN_X4M (D, GN, QN, SN);

	//ports
	input D;
	input GN;
	output QN;
	input SN;

	//wires
	wire D;
	wire GN;
	wire QN;
	wire SN;

endmodule


module LATQN_X0P5M (D, G, QN);

	//ports
	input D;
	input G;
	output QN;

	//wires
	wire D;
	wire G;
	wire QN;

endmodule


module LATQN_X1M (D, G, QN);

	//ports
	input D;
	input G;
	output QN;

	//wires
	wire D;
	wire G;
	wire QN;

endmodule


module LATQN_X2M (D, G, QN);

	//ports
	input D;
	input G;
	output QN;

	//wires
	wire D;
	wire G;
	wire QN;

endmodule


module LATQN_X3M (D, G, QN);

	//ports
	input D;
	input G;
	output QN;

	//wires
	wire D;
	wire G;
	wire QN;

endmodule


module LATQN_X4M (D, G, QN);

	//ports
	input D;
	input G;
	output QN;

	//wires
	wire D;
	wire G;
	wire QN;

endmodule


module LATQ_X0P5M (D, G, Q);

	//ports
	input D;
	input G;
	output Q;

	//wires
	wire D;
	wire G;
	wire Q;

endmodule


module LATQ_X1M (D, G, Q);

	//ports
	input D;
	input G;
	output Q;

	//wires
	wire D;
	wire G;
	wire Q;

endmodule


module LATQ_X2M (D, G, Q);

	//ports
	input D;
	input G;
	output Q;

	//wires
	wire D;
	wire G;
	wire Q;

endmodule


module LATQ_X3M (D, G, Q);

	//ports
	input D;
	input G;
	output Q;

	//wires
	wire D;
	wire G;
	wire Q;

endmodule


module LATRPQN_X0P5M (D, G, QN, R);

	//ports
	input D;
	input G;
	output QN;
	input R;

	//wires
	wire D;
	wire G;
	wire QN;
	wire R;

endmodule


module LATRPQN_X1M (D, G, QN, R);

	//ports
	input D;
	input G;
	output QN;
	input R;

	//wires
	wire D;
	wire G;
	wire QN;
	wire R;

endmodule


module LATRPQN_X2M (D, G, QN, R);

	//ports
	input D;
	input G;
	output QN;
	input R;

	//wires
	wire D;
	wire G;
	wire QN;
	wire R;

endmodule


module LATRPQN_X3M (D, G, QN, R);

	//ports
	input D;
	input G;
	output QN;
	input R;

	//wires
	wire D;
	wire G;
	wire QN;
	wire R;

endmodule


module LATRPQN_X4M (D, G, QN, R);

	//ports
	input D;
	input G;
	output QN;
	input R;

	//wires
	wire D;
	wire G;
	wire QN;
	wire R;

endmodule


module LATRQ_X0P5M (D, G, Q, RN);

	//ports
	input D;
	input G;
	output Q;
	input RN;

	//wires
	wire D;
	wire G;
	wire Q;
	wire RN;

endmodule


module LATRQ_X1M (D, G, Q, RN);

	//ports
	input D;
	input G;
	output Q;
	input RN;

	//wires
	wire D;
	wire G;
	wire Q;
	wire RN;

endmodule


module LATRQ_X2M (D, G, Q, RN);

	//ports
	input D;
	input G;
	output Q;
	input RN;

	//wires
	wire D;
	wire G;
	wire Q;
	wire RN;

endmodule


module LATRQ_X3M (D, G, Q, RN);

	//ports
	input D;
	input G;
	output Q;
	input RN;

	//wires
	wire D;
	wire G;
	wire Q;
	wire RN;

endmodule


module LATSPQ_X0P5M (D, G, Q, S);

	//ports
	input D;
	input G;
	output Q;
	input S;

	//wires
	wire D;
	wire G;
	wire Q;
	wire S;

endmodule


module LATSPQ_X1M (D, G, Q, S);

	//ports
	input D;
	input G;
	output Q;
	input S;

	//wires
	wire D;
	wire G;
	wire Q;
	wire S;

endmodule


module LATSPQ_X2M (D, G, Q, S);

	//ports
	input D;
	input G;
	output Q;
	input S;

	//wires
	wire D;
	wire G;
	wire Q;
	wire S;

endmodule


module LATSPQ_X3M (D, G, Q, S);

	//ports
	input D;
	input G;
	output Q;
	input S;

	//wires
	wire D;
	wire G;
	wire Q;
	wire S;

endmodule


module LATSQN_X0P5M (D, G, QN, SN);

	//ports
	input D;
	input G;
	output QN;
	input SN;

	//wires
	wire D;
	wire G;
	wire QN;
	wire SN;

endmodule


module LATSQN_X1M (D, G, QN, SN);

	//ports
	input D;
	input G;
	output QN;
	input SN;

	//wires
	wire D;
	wire G;
	wire QN;
	wire SN;

endmodule


module LATSQN_X2M (D, G, QN, SN);

	//ports
	input D;
	input G;
	output QN;
	input SN;

	//wires
	wire D;
	wire G;
	wire QN;
	wire SN;

endmodule


module LATSQN_X3M (D, G, QN, SN);

	//ports
	input D;
	input G;
	output QN;
	input SN;

	//wires
	wire D;
	wire G;
	wire QN;
	wire SN;

endmodule


module LATSQN_X4M (D, G, QN, SN);

	//ports
	input D;
	input G;
	output QN;
	input SN;

	//wires
	wire D;
	wire G;
	wire QN;
	wire SN;

endmodule


module M2DFFQN_X0P5M (CK, D0, D1, QN, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;

endmodule


module M2DFFQN_X1M (CK, D0, D1, QN, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;

endmodule


module M2DFFQN_X2M (CK, D0, D1, QN, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;

endmodule


module M2DFFQN_X3M (CK, D0, D1, QN, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;

endmodule


module M2DFFQ_X0P5M (CK, D0, D1, Q, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;

endmodule


module M2DFFQ_X1M (CK, D0, D1, Q, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;

endmodule


module M2DFFQ_X2M (CK, D0, D1, Q, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;

endmodule


module M2DFFQ_X3M (CK, D0, D1, Q, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;

endmodule


module M2DFFQ_X4M (CK, D0, D1, Q, S0);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;

endmodule


module M2SDFFQN_X0P5M (CK, D0, D1, QN, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQN_X1M (CK, D0, D1, QN, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQN_X2M (CK, D0, D1, QN, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQN_X3M (CK, D0, D1, QN, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output QN;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire QN;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQ_X0P5M (CK, D0, D1, Q, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQ_X1M (CK, D0, D1, Q, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQ_X2M (CK, D0, D1, Q, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQ_X3M (CK, D0, D1, Q, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;
	wire SE;
	wire SI;

endmodule


module M2SDFFQ_X4M (CK, D0, D1, Q, S0, SE, SI);

	//ports
	input CK;
	input D0;
	input D1;
	output Q;
	input S0;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D0;
	wire D1;
	wire Q;
	wire S0;
	wire SE;
	wire SI;

endmodule


module MX2_X0P5B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X0P5M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X0P7B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X0P7M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X1B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X1M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X1P4B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X1P4M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X2B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X2M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X3B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X3M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X4B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X4M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X6B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X6M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MX2_X8B (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X0P5M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X0P7M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X1M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X1P4M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X2M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X3M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT2_X4M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXIT4_X0P5M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXIT4_X0P7M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXIT4_X1M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXIT4_X1P4M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXIT4_X2M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXIT4_X3M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXT2_X0P5M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X0P7M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X1M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X1P4M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X2M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X3M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X4M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT2_X6M (A, B, S0, Y);

	//ports
	input A;
	input B;
	input S0;
	output Y;

	//wires
	wire A;
	wire B;
	wire S0;
	wire Y;

endmodule


module MXT4_X0P5M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXT4_X0P7M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXT4_X1M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXT4_X1P4M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXT4_X2M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module MXT4_X3M (A, B, C, D, S0, S1, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input S0;
	input S1;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire S0;
	wire S1;
	wire Y;

endmodule


module NAND2B_X0P5M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X0P7M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X1M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X1P4M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X2M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X3M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X4M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X6M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2B_X8M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NAND2XB_X0P5M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X0P7M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X1M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X1P4M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X2M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X3M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X4M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X6M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2XB_X8M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NAND2_X0P5A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X0P5B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X0P5M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X0P7A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X0P7B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X0P7M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X1A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X1B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X1M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X1P4A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X1P4B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X1P4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X2A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X2B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X2M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X3A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X3B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X3M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X4A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X4B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X6A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X6B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X6M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X8A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X8B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND2_X8M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NAND3B_X0P5M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X0P7M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X1M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X1P4M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X2M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X3M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X4M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3B_X6M (AN, B, C, Y);

	//ports
	input AN;
	input B;
	input C;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3XXB_X0P5M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X0P7M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X1M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X1P4M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X2M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X3M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X4M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3XXB_X6M (A, B, CN, Y);

	//ports
	input A;
	input B;
	input CN;
	output Y;

	//wires
	wire A;
	wire B;
	wire CN;
	wire Y;

endmodule


module NAND3_X0P5A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X0P5M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X0P7A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X0P7M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X1A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X1M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X1P4A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X1P4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X2A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X2M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X3A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X3M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X4A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X6A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND3_X6M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NAND4B_X0P5M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4B_X0P7M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4B_X1M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4B_X1P4M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4B_X2M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4B_X3M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4B_X4M (AN, B, C, D, Y);

	//ports
	input AN;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire AN;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4XXXB_X0P5M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4XXXB_X0P7M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4XXXB_X1M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4XXXB_X1P4M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4XXXB_X2M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4XXXB_X3M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4XXXB_X4M (A, B, C, DN, Y);

	//ports
	input A;
	input B;
	input C;
	input DN;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire DN;
	wire Y;

endmodule


module NAND4_X0P5A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X0P5M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X0P7A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X0P7M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X1A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X1M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X1P4A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X1P4M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X2A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X2M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X3A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X3M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X4A (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NAND4_X4M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module NOR2B_X0P5M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X0P7M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X1M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X1P4M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X2M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X3M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X4M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X6M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2B_X8M (AN, B, Y);

	//ports
	input AN;
	input B;
	output Y;

	//wires
	wire AN;
	wire B;
	wire Y;

endmodule


module NOR2XB_X0P5M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X0P7M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X1M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X1P4M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X2M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X3M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X4M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X6M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2XB_X8M (A, BN, Y);

	//ports
	input A;
	input BN;
	output Y;

	//wires
	wire A;
	wire BN;
	wire Y;

endmodule


module NOR2_X0P5A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X0P5B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X0P5M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X0P7A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X0P7B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X0P7M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X1A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X1B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X1M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X1P4A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X1P4B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X1P4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X2A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X2B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X2M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X3A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X3B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X3M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X4A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X4B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X6A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X6B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X6M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X8A (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X8B (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR2_X8M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module NOR3_X0P5A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X0P5M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X0P7A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X0P7M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X1A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X1M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X1P4A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X1P4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X2A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X2M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X3A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X3M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X4A (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module NOR3_X4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OA211_X0P5M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X0P7M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X1M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X1P4M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X2M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X3M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X4M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA211_X6M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OA21_X0P5M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X0P7M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X1M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X1P4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X2M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X3M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X6M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA21_X8M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OA22_X0P5M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X0P7M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X1M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X1P4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X2M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X3M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X6M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OA22_X8M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI211_X0P5M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI211_X0P7M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI211_X1M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI211_X1P4M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI211_X2M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI211_X3M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI211_X4M (A0, A1, B0, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire C0;
	wire Y;

endmodule


module OAI21B_X0P5M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X0P7M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X1M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X1P4M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X2M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X3M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X4M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X6M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21B_X8M (A0, A1, B0N, Y);

	//ports
	input A0;
	input A1;
	input B0N;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0N;
	wire Y;

endmodule


module OAI21_X0P5M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X0P7M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X1M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X1P4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X2M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X3M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X4M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X6M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI21_X8M (A0, A1, B0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire Y;

endmodule


module OAI221_X0P5M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI221_X0P7M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI221_X1M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI221_X1P4M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI221_X2M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI221_X3M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI221_X4M (A0, A1, B0, B1, C0, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire Y;

endmodule


module OAI222_X0P5M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI222_X0P7M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI222_X1M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI222_X1P4M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI222_X2M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI222_X3M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI222_X4M (A0, A1, B0, B1, C0, C1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	input C0;
	input C1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire C0;
	wire C1;
	wire Y;

endmodule


module OAI22_X0P5M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X0P7M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X1M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X1P4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X2M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X3M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X4M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X6M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI22_X8M (A0, A1, B0, B1, Y);

	//ports
	input A0;
	input A1;
	input B0;
	input B1;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire B0;
	wire B1;
	wire Y;

endmodule


module OAI2XB1_X0P5M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X0P7M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X1M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X1P4M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X2M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X3M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X4M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X6M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI2XB1_X8M (A0, A1N, B0, Y);

	//ports
	input A0;
	input A1N;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1N;
	wire B0;
	wire Y;

endmodule


module OAI31_X0P5M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X0P7M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X1M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X1P4M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X2M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X3M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X4M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OAI31_X6M (A0, A1, A2, B0, Y);

	//ports
	input A0;
	input A1;
	input A2;
	input B0;
	output Y;

	//wires
	wire A0;
	wire A1;
	wire A2;
	wire B0;
	wire Y;

endmodule


module OR2_X0P5M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X0P7M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X11M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X1M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X1P4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X2M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X3M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X6M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR2_X8M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module OR3_X0P5M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X0P7M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X1M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X1P4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X2M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X3M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X6M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR3_X8M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module OR4_X0P5M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X0P7M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X1M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X1P4M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X2M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X3M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X4M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X6M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR4_X8M (A, B, C, D, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire Y;

endmodule


module OR6_X0P5M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X0P7M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X1M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X1P4M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X2M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X3M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X4M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module OR6_X6M (A, B, C, D, E, F, Y);

	//ports
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire D;
	wire E;
	wire F;
	wire Y;

endmodule


module POSTICG_X0P5B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X0P6B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X0P7B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X0P8B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X11B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X13B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X16B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X1B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X1P2B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X1P4B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X1P7B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X2B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X2P5B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X3B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X3P5B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X4B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X5B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X6B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X7P5B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module POSTICG_X9B (CK, E, ECK, SEN);

	//ports
	input CK;
	input E;
	output ECK;
	input SEN;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SEN;

endmodule


module PREICG_X0P5B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X0P6B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X0P7B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X0P8B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X11B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X13B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X16B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X1B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X1P2B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X1P4B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X1P7B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X2B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X2P5B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X3B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X3P5B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X4B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X5B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X6B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X7P5B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module PREICG_X9B (CK, E, ECK, SE);

	//ports
	input CK;
	input E;
	output ECK;
	input SE;

	//wires
	wire CK;
	wire E;
	wire ECK;
	wire SE;

endmodule


module RF1R1WS_X1M (RBL, RWL, WBL, WWL);

	//ports
	output RBL;
	input RWL;
	input WBL;
	input WWL;

	//wires
	wire RBL;
	wire RWL;
	wire WBL;
	wire WWL;

endmodule


module RF1R1WS_X1P4M (RBL, RWL, WBL, WWL);

	//ports
	output RBL;
	input RWL;
	input WBL;
	input WWL;

	//wires
	wire RBL;
	wire RWL;
	wire WBL;
	wire WWL;

endmodule


module RF1R1WS_X2M (RBL, RWL, WBL, WWL);

	//ports
	output RBL;
	input RWL;
	input WBL;
	input WWL;

	//wires
	wire RBL;
	wire RWL;
	wire WBL;
	wire WWL;

endmodule


module RF1R2WS_X1M (RBL, RWL, WBL1, WBL2, WWL1, WWL2);

	//ports
	output RBL;
	input RWL;
	input WBL1;
	input WBL2;
	input WWL1;
	input WWL2;

	//wires
	wire RBL;
	wire RWL;
	wire WBL1;
	wire WBL2;
	wire WWL1;
	wire WWL2;

endmodule


module RF1R2WS_X1P4M (RBL, RWL, WBL1, WBL2, WWL1, WWL2);

	//ports
	output RBL;
	input RWL;
	input WBL1;
	input WBL2;
	input WWL1;
	input WWL2;

	//wires
	wire RBL;
	wire RWL;
	wire WBL1;
	wire WBL2;
	wire WWL1;
	wire WWL2;

endmodule


module RF1R2WS_X2M (RBL, RWL, WBL1, WBL2, WWL1, WWL2);

	//ports
	output RBL;
	input RWL;
	input WBL1;
	input WBL2;
	input WWL1;
	input WWL2;

	//wires
	wire RBL;
	wire RWL;
	wire WBL1;
	wire WBL2;
	wire WWL1;
	wire WWL2;

endmodule


module RF2R1WS_X1M (RBL1, RBL2, RWL1, RWL2, WBL, WWL);

	//ports
	output RBL1;
	output RBL2;
	input RWL1;
	input RWL2;
	input WBL;
	input WWL;

	//wires
	wire RBL1;
	wire RBL2;
	wire RWL1;
	wire RWL2;
	wire WBL;
	wire WWL;

endmodule


module RF2R1WS_X1P4M (RBL1, RBL2, RWL1, RWL2, WBL, WWL);

	//ports
	output RBL1;
	output RBL2;
	input RWL1;
	input RWL2;
	input WBL;
	input WWL;

	//wires
	wire RBL1;
	wire RBL2;
	wire RWL1;
	wire RWL2;
	wire WBL;
	wire WWL;

endmodule


module RF2R1WS_X2M (RBL1, RBL2, RWL1, RWL2, WBL, WWL);

	//ports
	output RBL1;
	output RBL2;
	input RWL1;
	input RWL2;
	input WBL;
	input WWL;

	//wires
	wire RBL1;
	wire RBL2;
	wire RWL1;
	wire RWL2;
	wire WBL;
	wire WWL;

endmodule


module RF2R2WS_X1M (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);

	//ports
	output RBL1;
	output RBL2;
	input RWL1;
	input RWL2;
	input WBL1;
	input WBL2;
	input WWL1;
	input WWL2;

	//wires
	wire RBL1;
	wire RBL2;
	wire RWL1;
	wire RWL2;
	wire WBL1;
	wire WBL2;
	wire WWL1;
	wire WWL2;

endmodule


module RF2R2WS_X1P4M (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);

	//ports
	output RBL1;
	output RBL2;
	input RWL1;
	input RWL2;
	input WBL1;
	input WBL2;
	input WWL1;
	input WWL2;

	//wires
	wire RBL1;
	wire RBL2;
	wire RWL1;
	wire RWL2;
	wire WBL1;
	wire WBL2;
	wire WWL1;
	wire WWL2;

endmodule


module RF2R2WS_X2M (RBL1, RBL2, RWL1, RWL2, WBL1, WBL2, WWL1, WWL2);

	//ports
	output RBL1;
	output RBL2;
	input RWL1;
	input RWL2;
	input WBL1;
	input WBL2;
	input WWL1;
	input WWL2;

	//wires
	wire RBL1;
	wire RBL2;
	wire RWL1;
	wire RWL2;
	wire WBL1;
	wire WBL2;
	wire WWL1;
	wire WWL2;

endmodule


module SDFFNQ_X1M (CKN, D, Q, SE, SI);

	//ports
	input CKN;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFNQ_X2M (CKN, D, Q, SE, SI);

	//ports
	input CKN;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFNQ_X3M (CKN, D, Q, SE, SI);

	//ports
	input CKN;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFNRPQ_X1M (CKN, D, Q, R, SE, SI);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFNRPQ_X2M (CKN, D, Q, R, SE, SI);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFNRPQ_X3M (CKN, D, Q, R, SE, SI);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFNSQ_X1M (CKN, D, Q, SE, SI, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFNSQ_X2M (CKN, D, Q, SE, SI, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFNSQ_X3M (CKN, D, Q, SE, SI, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFNSRPQ_X1M (CKN, D, Q, R, SE, SI, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFNSRPQ_X2M (CKN, D, Q, R, SE, SI, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFNSRPQ_X3M (CKN, D, Q, R, SE, SI, SN);

	//ports
	input CKN;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CKN;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFQN_X0P5M (CK, D, QN, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;

endmodule


module SDFFQN_X1M (CK, D, QN, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;

endmodule


module SDFFQN_X2M (CK, D, QN, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;

endmodule


module SDFFQN_X3M (CK, D, QN, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;

endmodule


module SDFFQ_X0P5M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFQ_X1M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFQ_X2M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFQ_X3M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFQ_X4M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFRPQN_X0P5M (CK, D, QN, R, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQN_X1M (CK, D, QN, R, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQN_X2M (CK, D, QN, R, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQN_X3M (CK, D, QN, R, SE, SI);

	//ports
	input CK;
	input D;
	output QN;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQ_X0P5M (CK, D, Q, R, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQ_X1M (CK, D, Q, R, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQ_X2M (CK, D, Q, R, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQ_X3M (CK, D, Q, R, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFRPQ_X4M (CK, D, Q, R, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;

endmodule


module SDFFSQN_X0P5M (CK, D, QN, SE, SI, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQN_X1M (CK, D, QN, SE, SI, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQN_X2M (CK, D, QN, SE, SI, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQN_X3M (CK, D, QN, SE, SI, SN);

	//ports
	input CK;
	input D;
	output QN;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire QN;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQ_X0P5M (CK, D, Q, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQ_X1M (CK, D, Q, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQ_X2M (CK, D, Q, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQ_X3M (CK, D, Q, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSQ_X4M (CK, D, Q, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSRPQ_X0P5M (CK, D, Q, R, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSRPQ_X1M (CK, D, Q, R, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSRPQ_X2M (CK, D, Q, R, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSRPQ_X3M (CK, D, Q, R, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFSRPQ_X4M (CK, D, Q, R, SE, SI, SN);

	//ports
	input CK;
	input D;
	output Q;
	input R;
	input SE;
	input SI;
	input SN;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire R;
	wire SE;
	wire SI;
	wire SN;

endmodule


module SDFFYQ_X1M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFYQ_X2M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFYQ_X3M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module SDFFYQ_X4M (CK, D, Q, SE, SI);

	//ports
	input CK;
	input D;
	output Q;
	input SE;
	input SI;

	//wires
	wire CK;
	wire D;
	wire Q;
	wire SE;
	wire SI;

endmodule


module TIEHI_X1M (Y);

	//ports
	output Y;

	//wires
	wire Y;

endmodule


module TIELO_X1M (Y);

	//ports
	output Y;

	//wires
	wire Y;

endmodule


module WELLANTENNATIEPW2 ();

	//wires

endmodule


module XNOR2_X0P5M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR2_X0P7M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR2_X1M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR2_X1P4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR2_X2M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR2_X3M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR2_X4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XNOR3_X0P5M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XNOR3_X0P7M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XNOR3_X1M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XNOR3_X1P4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XNOR3_X2M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XNOR3_X3M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XNOR3_X4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR2_X0P5M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR2_X0P7M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR2_X1M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR2_X1P4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR2_X2M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR2_X3M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR2_X4M (A, B, Y);

	//ports
	input A;
	input B;
	output Y;

	//wires
	wire A;
	wire B;
	wire Y;

endmodule


module XOR3_X0P5M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR3_X0P7M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR3_X1M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR3_X1P4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR3_X2M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR3_X3M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule


module XOR3_X4M (A, B, C, Y);

	//ports
	input A;
	input B;
	input C;
	output Y;

	//wires
	wire A;
	wire B;
	wire C;
	wire Y;

endmodule
